module and2
(
input in1_i,
input in2_i,

output reg out1_o
);

assign out1_o = in1_i & in2_i;

endmodule